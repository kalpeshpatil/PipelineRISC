library verilog;
use verilog.vl_types.all;
entity hazard_unit is
    port(
        IR_FD           : in     vl_logic_vector(15 downto 0);
        flush_FD        : out    vl_logic;
        flush_DR        : out    vl_logic;
        flush_RE        : out    vl_logic;
        flush_EM        : out    vl_logic;
        flush_MW        : out    vl_logic;
        flush_FD_in     : in     vl_logic;
        flush_DR_in     : in     vl_logic;
        flush_RE_in     : in     vl_logic;
        flush_EM_in     : in     vl_logic;
        flush_MW_in     : in     vl_logic;
        ALU_pc_muxA_ctrl: out    vl_logic;
        ALU_pc_muxB_ctrl: out    vl_logic;
        PC_mux_ctrl     : out    vl_logic_vector(2 downto 0);
        PC_en           : out    vl_logic;
        FD_en           : out    vl_logic;
        DR_en           : out    vl_logic;
        RE_en           : out    vl_logic;
        EM_en           : out    vl_logic;
        MW_en           : out    vl_logic;
        vbit_LM         : in     vl_logic;
        vbit_SM         : in     vl_logic;
        T3_ctrl         : out    vl_logic;
        R7_dest_RE      : in     vl_logic;
        R7_dest_EM      : in     vl_logic;
        R7_dest_MW      : in     vl_logic;
        load_RE         : in     vl_logic;
        load_EM         : in     vl_logic;
        load_MW         : in     vl_logic;
        LM_RE           : in     vl_logic;
        LM_EM           : in     vl_logic;
        LM_MW           : in     vl_logic;
        SM_DR           : in     vl_logic;
        SM_EM           : in     vl_logic;
        jump_bits_DR    : in     vl_logic_vector(1 downto 0);
        jump_bits_RE    : in     vl_logic_vector(1 downto 0);
        jump_bits_EM    : in     vl_logic_vector(1 downto 0);
        imm9FDctrl      : out    vl_logic;
        imm9EMctrl      : out    vl_logic;
        zero_flag       : in     vl_logic;
        store_RE        : in     vl_logic;
        reg_efct_RE     : in     vl_logic_vector(2 downto 0);
        reg_efct_EM     : in     vl_logic_vector(2 downto 0);
        Rd_MW           : in     vl_logic_vector(2 downto 0);
        Rd_EM           : in     vl_logic_vector(2 downto 0);
        Rs1_RE          : in     vl_logic_vector(2 downto 0);
        Rs2_RE          : in     vl_logic_vector(2 downto 0);
        prio_enc_LM_en  : out    vl_logic;
        prio_enc_SM_en  : out    vl_logic
    );
end hazard_unit;
