library verilog;
use verilog.vl_types.all;
entity se79_16 is
    port(
        \in\            : in     vl_logic_vector(8 downto 0);
        \out\           : out    vl_logic_vector(15 downto 0)
    );
end se79_16;
