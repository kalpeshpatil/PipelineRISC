library verilog;
use verilog.vl_types.all;
entity controller is
    port(
        clock           : in     vl_logic
    );
end controller;
